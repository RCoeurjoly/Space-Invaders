//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:30:38 03/19/2013 
// Design Name: 
// Module Name:    formatVGA
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module formatVGA(
		 input wire [9:0]  VGAx,
		 input wire [9:0]  VGAy,
		 input wire 	   clr, //asynchronous reset
		 input wire [19:0] invArray,
		 input wire [4:0]  invLine,
		 input wire [4:0]  shipX,
		 input wire [4:0]  bulletX,
		 input wire [3:0]  bulletY,
		 input wire 	   bulletFlying,
		 output reg [2:0]  rgb 
		 );   

   
   reg [31 : 0] 		   invader [31 : 0];
   reg [31 : 0] 		   ship [31 : 0];
   reg [31:0] 		   bullet [0:31];
   initial begin
      rgb <= 3'b000;
      
      invader[0] <= 32'b00000000000000000000000000000000;
      invader[1] <= 32'b00000000000000000000000000000000;
      invader[2] <= 32'b00000000000000000000000000000000;
      invader[3] <= 32'b00000000000000000000000000000000;
      invader[4] <= 32'b00000000000000000000000000000000;
      invader[5] <= 32'b00000000000000000000000000000000;
      invader[6] <= 32'b00000000000000000000000000000000;
      invader[7] <= 32'b00000000000000000000000000000000;
      invader[8] <= 32'b00000000011000000000011000000000;
      invader[9] <= 32'b00000000011000000000011000000000;
      invader[10] <= 32'b00000000000110000001100000000000;
      invader[11] <= 32'b00000000000110000001100000000000;
      invader[12] <= 32'b00000000011111111111111000000000;
      invader[13] <= 32'b00000000011111111111111000000000;
      invader[14] <= 32'b00000001111001111110011110000000;
      invader[15] <= 32'b00000001111001111110011110000000;
      invader[16] <= 32'b00000111111111111111111111100000;
      invader[17] <= 32'b00000111111111111111111111100000;
      invader[18] <= 32'b00000110011111111111111001100000;
      invader[19] <= 32'b00000110011111111111111001100000;
      invader[20] <= 32'b00000110011000000000011001100000;
      invader[21] <= 32'b00000110011000000000011001100000;
      invader[22] <= 32'b00000000000111100111100000000000;
      invader[23] <= 32'b00000000000111100111100000000000;
      invader[24] <= 32'b00000000000000000000000000000000;
      invader[25] <= 32'b00000000000000000000000000000000;
      invader[26] <= 32'b00000000000000000000000000000000;
      invader[27] <= 32'b00000000000000000000000000000000;
      invader[28] <= 32'b00000000000000000000000000000000;
      invader[29] <= 32'b00000000000000000000000000000000;
      invader[30] <= 32'b00000000000000000000000000000000;
      invader[31] <= 32'b00000000000000000000000000000000;
      
      ship[0] <= 32'b00000000000000011000000000000000;
      ship[1] <= 32'b00000000000000011000000000000000;
      ship[2] <= 32'b00000000000000011000000000000000;
      ship[3] <= 32'b00000000000000011000000000000000;
      ship[4] <= 32'b00000000000001111110000000000000;
      ship[5] <= 32'b00000000000001111110000000000000;
      ship[6] <= 32'b00000000000001111110000000000000;
      ship[7] <= 32'b00000000000001111110000000000000;
      ship[8] <= 32'b00000001100001111110000110000000;
      ship[9] <= 32'b00000001100001111110000110000000;
      ship[10] <= 32'b00000001100001111110000110000000;
      ship[11] <= 32'b00000001100001111110000110000000;
      ship[12] <= 32'b00000001100111111111100110000000;
      ship[13] <= 32'b00000001100111111111100110000000;
      ship[14] <= 32'b00000001111111100111111110000000;
      ship[15] <= 32'b00000001111111100111111110000000;
      ship[16] <= 32'b01100001111110000001111110000110;
      ship[17] <= 32'b01100001111110000001111110000110;
      ship[18] <= 32'b01100001111110000001111110000110;
      ship[19] <= 32'b01100001111110000001111110000110;
      ship[20] <= 32'b01100001111111111111111110000110;
      ship[21] <= 32'b01100001111111111111111110000110;
      ship[22] <= 32'b01100111111111111111111111100110;
      ship[23] <= 32'b01100111111111111111111111100110;
      ship[24] <= 32'b01111111111111111111111111111110;
      ship[25] <= 32'b01111111111111111111111111111110;
      ship[26] <= 32'b01111110011111111111111001111110;
      ship[27] <= 32'b01111110011111111111111001111110;
      ship[28] <= 32'b01111000011110011001111000011110;
      ship[29] <= 32'b01111000011110011001111000011110;
      ship[30] <= 32'b01100000000000011000000000000110;
      ship[31] <= 32'b01100000000000011000000000000110;

            
      bullet[0] <= 32'b00000000000000111100000000000000;
      bullet[1] <= 32'b00000000000001011110000000000000;
      bullet[2] <= 32'b00000000000010101111000000000000;
      bullet[3] <= 32'b00000000000110001111100000000000;
      bullet[4] <= 32'b00000000001111111111110000000000;
      bullet[5] <= 32'b00000000001111110011110000000000;
      bullet[6] <= 32'b00000000011111110001111000000000;
      bullet[7] <= 32'b00000000011111100001111000000000;
      bullet[8] <= 32'b00000000011111110001111000000000;
      bullet[9] <= 32'b00000000011111100001111000000000;
      bullet[10] <= 32'b00000000011111100011111000000000;
      bullet[11] <= 32'b00000000011111110011111000000000;
      bullet[12] <= 32'b00000000011111111111111000000000;
      bullet[13] <= 32'b00000000000000000000000000000000;
      bullet[14] <= 32'b00000000010111111111111000000000;
      bullet[15] <= 32'b00000000010111111111111000000000;
      bullet[16] <= 32'b00000000000000000000000000000000;
      bullet[17] <= 32'b00000000000000000000000000000000;
      bullet[18] <= 32'b00000000000000000000000000000000;
      bullet[19] <= 32'b00000000000000000000000000000000;
      bullet[20] <= 32'b00000000000000000000000000000000;
      bullet[21] <= 32'b00000000000000000000000000000000;
      bullet[22] <= 32'b00000000000000000000000000000000;
      bullet[23] <= 32'b00000000000000000000000000000000;
      bullet[24] <= 32'b00000000000000000000000000000000;
      bullet[25] <= 32'b00000000000000000000000000000000;
      bullet[26] <= 32'b00000000000000000000000000000000;
      bullet[27] <= 32'b00000000000000000000000000000000;
      bullet[28] <= 32'b00000000000000000000000000000000;
      bullet[29] <= 32'b00000000000000000000000000000000;
      bullet[30] <= 32'b00000000000000000000000000000000;
      bullet[31] <= 32'b00000000000000000000000000000000;
      /**/
   end
   
   parameter [2:0] 	   black = 3'b000;
   parameter [2:0] 	   blue = 3'b001;
   parameter [2:0] 	   green = 3'b010;
   parameter [2:0] 	   cyan = 3'b011;
   parameter [2:0] 	   red = 3'b100;
   parameter [2:0] 	   magenta = 3'b101;
   parameter [2:0] 	   yellow = 3'b110;
   parameter [2:0] 	   white = 3'b111;
   
   wire [4:0] 			   x = VGAx[9:5];
   wire [3:0] 			   y = VGAy[8:5];
   wire [4:0] 			   indX = VGAx[4:0];
   wire [4:0] 			   indY = VGAy[4:0];
   reg [5:0] 			   indInv;
   reg [1:0] 			   currentInvader;
   reg 				   currentPixel;
   
   always @(*)
     begin
	if (clr == 1)
	  begin
	     // drawing bullet
	     if (bulletFlying == 1 && (x == bulletX) && (y == bulletY))
	       begin
		  if (bullet[indY][indX] == 1)
		    rgb <= yellow;
		  else
		    rgb <= black;
	       end
	     // drawing ship
	     else if (x == shipX && y == 13)
	       begin
		  if (ship[indY][indX] == 1)
		    rgb <= red;
		  else
		    rgb <= black;
	       end
	     // drawing invader
	     else if (y == invLine && invArray[x] == 1)
	       begin
		  if (invader[indY][indX] == 1)
		    rgb <= magenta;
		  else
		    rgb <= black;
	       end
	     //background
	     else
	       rgb <= black;/**/
	  end // if (clr == 1)
	else 
	  begin 
	     if (x[0] ^ y[0] == 1)
	       rgb <= white;
	     else rgb <= black;
	  end
     end // always @ (*)
   
   
   //end
endmodule
